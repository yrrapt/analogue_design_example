**.subckt auto_dac_unit_cell_test
**.ends
** flattened .save nodes
.end
